`ifdef ALU_LOADED
`else
`define ALU_LOADED

`include "./ALU/Add.sv"
`include "./ALU/Sub.sv"

`endif
